##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Sun May 29 22:07:47 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO user_proj_example
  CLASS BLOCK ;
  SIZE 823.860000 BY 814.640000 ;
  FOREIGN user_proj_example 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.852 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.57 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 86.7636 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 463.68 LAYER met3  ;
    ANTENNAGATEAREA 0.852 LAYER met3  ;
    ANTENNAMAXAREACAR 102.795 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 547.98 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.107277 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1.615000 0.000000 1.755000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.408 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 19.0413 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.4643 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.620000 0.000000 0.760000 0.490000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.065000 0.000000 175.205000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.870000 0.000000 59.010000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.750000 0.000000 176.890000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.380000 0.000000 173.520000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.700000 0.000000 171.840000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.015000 0.000000 170.155000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.330000 0.000000 168.470000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.760000 0.000000 112.900000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.075000 0.000000 111.215000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.390000 0.000000 109.530000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.705000 0.000000 107.845000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.020000 0.000000 106.160000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.340000 0.000000 104.480000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.655000 0.000000 102.795000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.970000 0.000000 101.110000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.285000 0.000000 99.425000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.600000 0.000000 97.740000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.920000 0.000000 96.060000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.235000 0.000000 94.375000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550000 0.000000 92.690000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.865000 0.000000 91.005000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.180000 0.000000 89.320000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.500000 0.000000 87.640000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.815000 0.000000 85.955000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.130000 0.000000 84.270000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.445000 0.000000 82.585000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.760000 0.000000 80.900000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.080000 0.000000 79.220000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.395000 0.000000 77.535000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.710000 0.000000 75.850000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.025000 0.000000 74.165000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.340000 0.000000 72.480000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.660000 0.000000 70.800000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.975000 0.000000 69.115000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.290000 0.000000 67.430000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.605000 0.000000 65.745000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.920000 0.000000 64.060000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.240000 0.000000 62.380000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.555000 0.000000 60.695000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.185000 0.000000 57.325000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.500000 0.000000 55.640000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.820000 0.000000 53.960000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.135000 0.000000 52.275000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.450000 0.000000 50.590000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.765000 0.000000 48.905000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.080000 0.000000 47.220000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.400000 0.000000 45.540000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.715000 0.000000 43.855000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.030000 0.000000 42.170000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.345000 0.000000 40.485000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.660000 0.000000 38.800000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.980000 0.000000 37.120000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.295000 0.000000 35.435000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.610000 0.000000 33.750000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.925000 0.000000 32.065000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.240000 0.000000 30.380000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.560000 0.000000 28.700000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.875000 0.000000 27.015000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.190000 0.000000 25.330000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.505000 0.000000 23.645000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.820000 0.000000 21.960000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.140000 0.000000 20.280000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.455000 0.000000 18.595000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.770000 0.000000 16.910000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.085000 0.000000 15.225000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.400000 0.000000 13.540000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.720000 0.000000 11.860000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.035000 0.000000 10.175000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.350000 0.000000 8.490000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.665000 0.000000 6.805000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.980000 0.000000 5.120000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 3.300000 0.000000 3.440000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 166.645000 0.000000 166.785000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 164.960000 0.000000 165.100000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 163.280000 0.000000 163.420000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 161.595000 0.000000 161.735000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 159.910000 0.000000 160.050000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 158.225000 0.000000 158.365000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 156.540000 0.000000 156.680000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 154.860000 0.000000 155.000000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 153.175000 0.000000 153.315000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 151.490000 0.000000 151.630000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 149.805000 0.000000 149.945000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 148.120000 0.000000 148.260000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 146.440000 0.000000 146.580000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 144.755000 0.000000 144.895000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 143.070000 0.000000 143.210000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 141.385000 0.000000 141.525000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 139.700000 0.000000 139.840000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 138.020000 0.000000 138.160000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 136.335000 0.000000 136.475000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 134.650000 0.000000 134.790000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 132.965000 0.000000 133.105000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 131.280000 0.000000 131.420000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 129.600000 0.000000 129.740000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 127.915000 0.000000 128.055000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 126.230000 0.000000 126.370000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 124.545000 0.000000 124.685000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 122.860000 0.000000 123.000000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 121.180000 0.000000 121.320000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 119.495000 0.000000 119.635000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 117.810000 0.000000 117.950000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 116.125000 0.000000 116.265000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.3025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 114.440000 0.000000 114.580000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.300000 0.000000 392.440000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.620000 0.000000 390.760000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.935000 0.000000 389.075000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.250000 0.000000 387.390000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.565000 0.000000 385.705000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.880000 0.000000 384.020000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.200000 0.000000 382.340000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.515000 0.000000 380.655000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.830000 0.000000 378.970000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.145000 0.000000 377.285000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.460000 0.000000 375.600000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.780000 0.000000 373.920000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.095000 0.000000 372.235000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.410000 0.000000 370.550000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.725000 0.000000 368.865000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.040000 0.000000 367.180000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.360000 0.000000 365.500000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.675000 0.000000 363.815000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.990000 0.000000 362.130000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.305000 0.000000 360.445000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.620000 0.000000 358.760000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.940000 0.000000 357.080000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.255000 0.000000 355.395000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.570000 0.000000 353.710000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.885000 0.000000 352.025000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.200000 0.000000 350.340000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.520000 0.000000 348.660000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.835000 0.000000 346.975000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.150000 0.000000 345.290000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.465000 0.000000 343.605000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.780000 0.000000 341.920000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.100000 0.000000 340.240000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.415000 0.000000 338.555000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.730000 0.000000 336.870000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.045000 0.000000 335.185000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.360000 0.000000 333.500000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.680000 0.000000 331.820000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.995000 0.000000 330.135000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.310000 0.000000 328.450000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.625000 0.000000 326.765000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.940000 0.000000 325.080000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.260000 0.000000 323.400000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.575000 0.000000 321.715000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.890000 0.000000 320.030000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.205000 0.000000 318.345000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.520000 0.000000 316.660000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.840000 0.000000 314.980000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.155000 0.000000 313.295000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.470000 0.000000 311.610000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.785000 0.000000 309.925000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.100000 0.000000 308.240000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.420000 0.000000 306.560000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.735000 0.000000 304.875000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.050000 0.000000 303.190000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.365000 0.000000 301.505000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.680000 0.000000 299.820000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.000000 0.000000 298.140000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.315000 0.000000 296.455000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.630000 0.000000 294.770000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.945000 0.000000 293.085000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.260000 0.000000 291.400000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.580000 0.000000 289.720000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5715 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 2.28737 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.84748 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0519192 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 287.895000 0.000000 288.035000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 342.967 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1839.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 10.5795 LAYER met4  ;
    ANTENNAMAXAREACAR 106.158 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 563.799 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.692525 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 286.210000 0.000000 286.350000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.525000 0.000000 284.665000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.840000 0.000000 282.980000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.160000 0.000000 281.300000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.475000 0.000000 279.615000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.790000 0.000000 277.930000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.105000 0.000000 276.245000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.420000 0.000000 274.560000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.740000 0.000000 272.880000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.055000 0.000000 271.195000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.370000 0.000000 269.510000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.685000 0.000000 267.825000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.000000 0.000000 266.140000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.320000 0.000000 264.460000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.635000 0.000000 262.775000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.950000 0.000000 261.090000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.265000 0.000000 259.405000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.580000 0.000000 257.720000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.900000 0.000000 256.040000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.215000 0.000000 254.355000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.530000 0.000000 252.670000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.845000 0.000000 250.985000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.160000 0.000000 249.300000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.480000 0.000000 247.620000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.795000 0.000000 245.935000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.110000 0.000000 244.250000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.425000 0.000000 242.565000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.740000 0.000000 240.880000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.060000 0.000000 239.200000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.375000 0.000000 237.515000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.690000 0.000000 235.830000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.005000 0.000000 234.145000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.320000 0.000000 232.460000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.640000 0.000000 230.780000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.955000 0.000000 229.095000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.270000 0.000000 227.410000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.585000 0.000000 225.725000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.900000 0.000000 224.040000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.220000 0.000000 222.360000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.535000 0.000000 220.675000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.850000 0.000000 218.990000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.165000 0.000000 217.305000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.480000 0.000000 215.620000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.800000 0.000000 213.940000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.115000 0.000000 212.255000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.430000 0.000000 210.570000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.745000 0.000000 208.885000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.060000 0.000000 207.200000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.380000 0.000000 205.520000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.695000 0.000000 203.835000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.010000 0.000000 202.150000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.325000 0.000000 200.465000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.640000 0.000000 198.780000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.960000 0.000000 197.100000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.275000 0.000000 195.415000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.590000 0.000000 193.730000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.905000 0.000000 192.045000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.220000 0.000000 190.360000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.540000 0.000000 188.680000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.855000 0.000000 186.995000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.170000 0.000000 185.310000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.485000 0.000000 183.625000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.800000 0.000000 181.940000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7798 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.673 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.6261 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.9969 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 180.120000 0.000000 180.260000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.435000 0.000000 178.575000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.6944 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.291 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 607.855000 0.000000 607.995000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 606.170000 0.000000 606.310000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 604.485000 0.000000 604.625000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 602.800000 0.000000 602.940000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 601.120000 0.000000 601.260000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 599.435000 0.000000 599.575000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 597.750000 0.000000 597.890000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 596.065000 0.000000 596.205000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 594.380000 0.000000 594.520000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 592.700000 0.000000 592.840000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 591.015000 0.000000 591.155000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 589.330000 0.000000 589.470000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 587.645000 0.000000 587.785000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 585.960000 0.000000 586.100000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 584.280000 0.000000 584.420000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 582.595000 0.000000 582.735000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 580.910000 0.000000 581.050000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 579.225000 0.000000 579.365000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 577.540000 0.000000 577.680000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 575.860000 0.000000 576.000000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 574.175000 0.000000 574.315000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 572.490000 0.000000 572.630000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 570.805000 0.000000 570.945000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 569.120000 0.000000 569.260000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 567.440000 0.000000 567.580000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 565.755000 0.000000 565.895000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 564.070000 0.000000 564.210000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 562.385000 0.000000 562.525000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 560.700000 0.000000 560.840000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 559.020000 0.000000 559.160000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 557.335000 0.000000 557.475000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 555.650000 0.000000 555.790000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 553.965000 0.000000 554.105000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 552.280000 0.000000 552.420000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 550.600000 0.000000 550.740000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 548.915000 0.000000 549.055000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 547.230000 0.000000 547.370000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 545.545000 0.000000 545.685000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 543.860000 0.000000 544.000000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 542.180000 0.000000 542.320000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 540.495000 0.000000 540.635000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 538.810000 0.000000 538.950000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 537.125000 0.000000 537.265000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 535.440000 0.000000 535.580000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 533.760000 0.000000 533.900000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 532.075000 0.000000 532.215000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 530.390000 0.000000 530.530000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 528.705000 0.000000 528.845000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 527.020000 0.000000 527.160000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 525.340000 0.000000 525.480000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 523.655000 0.000000 523.795000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 521.970000 0.000000 522.110000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 520.285000 0.000000 520.425000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 518.600000 0.000000 518.740000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 516.920000 0.000000 517.060000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 515.235000 0.000000 515.375000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 513.550000 0.000000 513.690000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 511.865000 0.000000 512.005000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 510.180000 0.000000 510.320000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 508.500000 0.000000 508.640000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 506.815000 0.000000 506.955000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 505.130000 0.000000 505.270000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 503.445000 0.000000 503.585000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 501.760000 0.000000 501.900000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 500.080000 0.000000 500.220000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 498.395000 0.000000 498.535000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 496.710000 0.000000 496.850000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 495.025000 0.000000 495.165000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 493.340000 0.000000 493.480000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 491.660000 0.000000 491.800000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 489.975000 0.000000 490.115000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 488.290000 0.000000 488.430000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 486.605000 0.000000 486.745000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 484.920000 0.000000 485.060000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 483.240000 0.000000 483.380000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 481.555000 0.000000 481.695000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 479.870000 0.000000 480.010000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 478.185000 0.000000 478.325000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 476.500000 0.000000 476.640000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 474.820000 0.000000 474.960000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 473.135000 0.000000 473.275000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 471.450000 0.000000 471.590000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 469.765000 0.000000 469.905000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 468.080000 0.000000 468.220000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 466.400000 0.000000 466.540000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 464.715000 0.000000 464.855000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 463.030000 0.000000 463.170000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 461.345000 0.000000 461.485000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 459.660000 0.000000 459.800000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 457.980000 0.000000 458.120000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 456.295000 0.000000 456.435000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 454.610000 0.000000 454.750000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 452.925000 0.000000 453.065000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 451.240000 0.000000 451.380000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 449.560000 0.000000 449.700000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.6944 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.291 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 447.875000 0.000000 448.015000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7329 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.3348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 290.256 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 446.190000 0.000000 446.330000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2812 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.4198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 285.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 444.505000 0.000000 444.645000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.1011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.3445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.3788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 231.824 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 442.820000 0.000000 442.960000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7147 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.2628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 305.872 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 441.140000 0.000000 441.280000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0274 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.976 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.3918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 242.56 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 439.455000 0.000000 439.595000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.3625 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.6515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.01 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.7668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 196.56 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 437.770000 0.000000 437.910000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.43 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.091 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.3898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 221.216 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 436.085000 0.000000 436.225000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.3828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 290.512 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 434.400000 0.000000 434.540000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8349 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.0135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.714 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.1368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 241.2 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 432.720000 0.000000 432.860000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.733 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.7928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 218.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 431.035000 0.000000 431.175000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4238 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.958 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.2608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 284.528 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 429.350000 0.000000 429.490000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2919 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.286 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 62.4588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 333.584 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 427.665000 0.000000 427.805000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4179 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.9285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.772 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.1478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 246.592 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 425.980000 0.000000 426.120000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8531 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.1045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.0408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 272.688 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 424.300000 0.000000 424.440000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.866 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.542 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.2108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 294.928 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 422.615000 0.000000 422.755000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1265 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.4715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.3568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 269.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 420.930000 0.000000 421.070000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 419.245000 0.000000 419.385000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 417.560000 0.000000 417.700000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 415.880000 0.000000 416.020000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 414.195000 0.000000 414.335000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 412.510000 0.000000 412.650000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 410.825000 0.000000 410.965000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 409.140000 0.000000 409.280000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 407.460000 0.000000 407.600000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 405.775000 0.000000 405.915000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 404.090000 0.000000 404.230000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 402.405000 0.000000 402.545000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 400.720000 0.000000 400.860000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 399.040000 0.000000 399.180000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.393 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 397.355000 0.000000 397.495000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 395.670000 0.000000 395.810000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.6846 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.144 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 393.985000 0.000000 394.125000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.180000 0.000000 822.320000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.720000 0.000000 821.860000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.040000 0.000000 820.180000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.355000 0.000000 818.495000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.670000 0.000000 816.810000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.985000 0.000000 815.125000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.300000 0.000000 813.440000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.620000 0.000000 811.760000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.935000 0.000000 810.075000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.250000 0.000000 808.390000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.565000 0.000000 806.705000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.880000 0.000000 805.020000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.200000 0.000000 803.340000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.515000 0.000000 801.655000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.830000 0.000000 799.970000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.145000 0.000000 798.285000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.460000 0.000000 796.600000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.780000 0.000000 794.920000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.095000 0.000000 793.235000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.410000 0.000000 791.550000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.725000 0.000000 789.865000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.040000 0.000000 788.180000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.360000 0.000000 786.500000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.675000 0.000000 784.815000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.990000 0.000000 783.130000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.305000 0.000000 781.445000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.620000 0.000000 779.760000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.940000 0.000000 778.080000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.255000 0.000000 776.395000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.570000 0.000000 774.710000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.885000 0.000000 773.025000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.200000 0.000000 771.340000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.520000 0.000000 769.660000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.835000 0.000000 767.975000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.150000 0.000000 766.290000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.465000 0.000000 764.605000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.780000 0.000000 762.920000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.100000 0.000000 761.240000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.415000 0.000000 759.555000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.730000 0.000000 757.870000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.045000 0.000000 756.185000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.360000 0.000000 754.500000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.680000 0.000000 752.820000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.995000 0.000000 751.135000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.310000 0.000000 749.450000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.625000 0.000000 747.765000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.940000 0.000000 746.080000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.260000 0.000000 744.400000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.575000 0.000000 742.715000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.890000 0.000000 741.030000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.205000 0.000000 739.345000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.520000 0.000000 737.660000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.840000 0.000000 735.980000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.155000 0.000000 734.295000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.470000 0.000000 732.610000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.785000 0.000000 730.925000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.100000 0.000000 729.240000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.420000 0.000000 727.560000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.735000 0.000000 725.875000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.050000 0.000000 724.190000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.365000 0.000000 722.505000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.680000 0.000000 720.820000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2106 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.591 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 9.32222 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.6596 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.162222 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 719.000000 0.000000 719.140000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.481 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 205.553 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1101.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 16.0245 LAYER met4  ;
    ANTENNAMAXAREACAR 40.272 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 209.545 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.340391 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 717.315000 0.000000 717.455000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.630000 0.000000 715.770000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.945000 0.000000 714.085000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.260000 0.000000 712.400000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.580000 0.000000 710.720000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.895000 0.000000 709.035000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.210000 0.000000 707.350000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.525000 0.000000 705.665000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.840000 0.000000 703.980000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.160000 0.000000 702.300000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.475000 0.000000 700.615000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.790000 0.000000 698.930000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.105000 0.000000 697.245000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.420000 0.000000 695.560000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.740000 0.000000 693.880000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.055000 0.000000 692.195000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.370000 0.000000 690.510000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.685000 0.000000 688.825000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.000000 0.000000 687.140000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.320000 0.000000 685.460000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.635000 0.000000 683.775000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.950000 0.000000 682.090000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.265000 0.000000 680.405000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.580000 0.000000 678.720000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.900000 0.000000 677.040000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.215000 0.000000 675.355000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530000 0.000000 673.670000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.845000 0.000000 671.985000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.160000 0.000000 670.300000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.480000 0.000000 668.620000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.795000 0.000000 666.935000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.110000 0.000000 665.250000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.425000 0.000000 663.565000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.826 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.85172 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.996 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 661.740000 0.000000 661.880000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.722 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.64566 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.1919 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 660.060000 0.000000 660.200000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6195 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.59717 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.9313 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 658.375000 0.000000 658.515000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.547 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.05788 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.1232 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 656.690000 0.000000 656.830000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.826 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.68485 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.1616 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 655.005000 0.000000 655.145000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7884 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.834 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.47596 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.3434 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 653.320000 0.000000 653.460000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.015 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.39636 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.9273 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 651.640000 0.000000 651.780000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.52 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.84414 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.0545 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 649.955000 0.000000 650.095000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6946 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.365 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.1899 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.6869 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 648.270000 0.000000 648.410000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7471 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6275 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.84727 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.4727 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 646.585000 0.000000 646.725000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.714 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 7.95152 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.9758 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 644.900000 0.000000 645.040000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6848 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.316 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.91202 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.3939 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 643.220000 0.000000 643.360000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5015 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.82061 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.8404 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 641.535000 0.000000 641.675000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7702 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.743 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.40242 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.9758 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 639.850000 0.000000 639.990000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3755 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 7.72707 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.7556 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 638.165000 0.000000 638.305000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7268 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.526 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.30111 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.3394 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 636.480000 0.000000 636.620000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.800000 0.000000 634.940000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.115000 0.000000 633.255000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.430000 0.000000 631.570000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.745000 0.000000 629.885000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.060000 0.000000 628.200000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.380000 0.000000 626.520000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.695000 0.000000 624.835000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.010000 0.000000 623.150000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.325000 0.000000 621.465000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.640000 0.000000 619.780000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.960000 0.000000 618.100000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.275000 0.000000 616.415000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.590000 0.000000 614.730000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.905000 0.000000 613.045000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.826 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 8.60283 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.4984 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.161635 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 611.220000 0.000000 611.360000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.540000 0.000000 609.680000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 39.590000 0.800000 39.890000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 99.195000 0.800000 99.495000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 158.800000 0.800000 159.100000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 218.410000 0.800000 218.710000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 278.015000 0.800000 278.315000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 337.625000 0.800000 337.925000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 397.230000 0.800000 397.530000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 456.835000 0.800000 457.135000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 516.445000 0.800000 516.745000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 576.050000 0.800000 576.350000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 635.660000 0.800000 635.960000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 695.265000 0.800000 695.565000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 754.870000 0.800000 755.170000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 810.540000 0.800000 810.840000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.300000 814.150000 63.440000 814.640000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.360000 814.150000 158.500000 814.640000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.420000 814.150000 253.560000 814.640000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.475000 814.150000 348.615000 814.640000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.535000 814.150000 443.675000 814.640000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.590000 814.150000 538.730000 814.640000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.650000 814.150000 633.790000 814.640000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.710000 814.150000 728.850000 814.640000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.800000 814.150000 820.940000 814.640000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.060000 777.440000 823.860000 777.740000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.060000 721.895000 823.860000 722.195000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.060000 666.355000 823.860000 666.655000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.060000 610.810000 823.860000 611.110000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.060000 555.270000 823.860000 555.570000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.060000 499.730000 823.860000 500.030000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.060000 444.185000 823.860000 444.485000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.060000 388.645000 823.860000 388.945000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.060000 333.100000 823.860000 333.400000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.8414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 271.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 47.4277 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 243.736 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 277.560000 823.860000 277.860000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.060000 222.020000 823.860000 222.320000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.060000 166.475000 823.860000 166.775000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.060000 110.935000 823.860000 111.235000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.060000 55.390000 823.860000 55.690000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.060000 9.610000 823.860000 9.910000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4923 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 19.720000 0.800000 20.020000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 79.325000 0.800000 79.625000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8641 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 138.935000 0.800000 139.235000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9136 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 198.540000 0.800000 198.840000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7591 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 258.145000 0.800000 258.445000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0171 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 317.755000 0.800000 318.055000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 377.360000 0.800000 377.660000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 436.970000 0.800000 437.270000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 496.575000 0.800000 496.875000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 556.180000 0.800000 556.480000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 615.790000 0.800000 616.090000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 675.395000 0.800000 675.695000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 735.005000 0.800000 735.305000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 794.610000 0.800000 794.910000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.628 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.979 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 54.634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 291.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 156.221 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 833.648 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 31.615000 814.150000 31.755000 814.640000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.5616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 122.647 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.616 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 125.578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 670.688 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 126.675000 814.150000 126.815000 814.640000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.9049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.364 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 123.479 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 659.024 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 221.730000 814.150000 221.870000 814.640000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7539 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 178.624 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 953.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 316.790000 814.150000 316.930000 814.640000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1372 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 34.945 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 186.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 175.004 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 933.824 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 411.850000 814.150000 411.990000 814.640000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.62 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.664 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.7396 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 223.552 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 506.905000 814.150000 507.045000 814.640000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.5365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.06 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.3918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 226.56 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 601.965000 814.150000 602.105000 814.640000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.452 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.7318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 207.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 697.020000 814.150000 697.160000 814.640000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7609 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 165.766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 885.024 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 792.080000 814.150000 792.220000 814.640000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 104.58 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 558.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.9958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 208.448 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 795.950000 823.860000 796.250000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 109.587 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 584.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.3418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 252.96 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 740.410000 823.860000 740.710000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.8304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.6668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 153.36 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 684.870000 823.860000 685.170000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5289 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.9238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 176.064 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 629.325000 823.860000 629.625000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4789 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.9518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 234.88 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 573.785000 823.860000 574.085000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.9408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 229.488 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 518.240000 823.860000 518.540000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 107.142 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 571.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.5398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 254.016 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 462.700000 823.860000 463.000000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 407.160000 823.860000 407.460000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 351.615000 823.860000 351.915000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 296.075000 823.860000 296.375000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 240.530000 823.860000 240.830000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 184.990000 823.860000 185.290000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 129.450000 823.860000 129.750000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 73.905000 823.860000 74.205000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 18.365000 823.860000 18.665000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4473 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 10.220000 0.800000 10.520000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 59.455000 0.800000 59.755000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9661 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 119.065000 0.800000 119.365000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 178.670000 0.800000 178.970000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1206 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 238.280000 0.800000 238.580000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7861 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 297.885000 0.800000 298.185000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.611 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1222.5 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 357.490000 0.800000 357.790000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 417.100000 0.800000 417.400000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 476.705000 0.800000 477.005000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 536.315000 0.800000 536.615000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 595.920000 0.800000 596.220000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 655.525000 0.800000 655.825000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 715.135000 0.800000 715.435000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 774.740000 0.800000 775.040000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.532 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 10.280000 814.150000 10.420000 814.640000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1288 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.483 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 94.990000 814.150000 95.130000 814.640000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 190.045000 814.150000 190.185000 814.640000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 285.105000 814.150000 285.245000 814.640000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 380.160000 814.150000 380.300000 814.640000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 475.220000 814.150000 475.360000 814.640000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 570.280000 814.150000 570.420000 814.640000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 665.335000 814.150000 665.475000 814.640000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.148 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 760.395000 814.150000 760.535000 814.640000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.641 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1222.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 809.930000 823.860000 810.230000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 758.925000 823.860000 759.225000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 703.380000 823.860000 703.680000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 647.840000 823.860000 648.140000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 592.300000 823.860000 592.600000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 536.755000 823.860000 537.055000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 481.215000 823.860000 481.515000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 425.670000 823.860000 425.970000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 370.130000 823.860000 370.430000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 69.1751 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 370.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.654 LAYER met4  ;
    ANTENNAMAXAREACAR 90.9071 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 475.636 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 314.590000 823.860000 314.890000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 259.045000 823.860000 259.345000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 203.505000 823.860000 203.805000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 147.960000 823.860000 148.260000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 92.420000 823.860000 92.720000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1221.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 823.060000 36.880000 823.860000 37.180000 ;
    END
  END io_oeb[0]
  PIN irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0048 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 322.385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.68 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1.080000 814.155000 1.220000 814.640000 ;
    END
  END irq[2]
  PIN irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0048 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 322.385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.68 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.620000 814.155000 0.760000 814.640000 ;
    END
  END irq[1]
  PIN irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 64.9852 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 322.189 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.68 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 225.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1223.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 105.971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.160000 814.155000 0.300000 814.640000 ;
    END
  END irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 815.800000 6.100000 817.800000 808.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.800000 0.800000 817.000000 6.100000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.060000 6.100000 8.060000 808.540000 ;
    END
    PORT
      LAYER met3 ;
        RECT 821.860000 382.450000 823.860000 384.450000 ;
    END
    PORT
      LAYER met4 ;
        RECT 309.465000 812.640000 311.465000 814.640000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 789.145000 386.810000 790.885000 781.590000 ;
      LAYER met4 ;
        RECT 313.825000 386.810000 315.565000 781.590000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 819.800000 2.100000 821.800000 812.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.060000 2.100000 4.060000 812.540000 ;
    END
    PORT
      LAYER met3 ;
        RECT 821.860000 378.450000 823.860000 380.450000 ;
    END
    PORT
      LAYER met4 ;
        RECT 305.465000 812.640000 307.465000 814.640000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 317.225000 390.210000 318.965000 778.190000 ;
      LAYER met4 ;
        RECT 785.745000 390.210000 787.485000 778.190000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 823.860000 814.640000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 823.860000 814.640000 ;
    LAYER met2 ;
      RECT 1.360000 814.015000 10.140000 814.640000 ;
      RECT 0.900000 814.015000 0.940000 814.640000 ;
      RECT 0.440000 814.015000 0.480000 814.640000 ;
      RECT 0.000000 814.015000 0.020000 814.640000 ;
      RECT 821.080000 814.010000 823.860000 814.640000 ;
      RECT 792.360000 814.010000 820.660000 814.640000 ;
      RECT 760.675000 814.010000 791.940000 814.640000 ;
      RECT 728.990000 814.010000 760.255000 814.640000 ;
      RECT 697.300000 814.010000 728.570000 814.640000 ;
      RECT 665.615000 814.010000 696.880000 814.640000 ;
      RECT 633.930000 814.010000 665.195000 814.640000 ;
      RECT 602.245000 814.010000 633.510000 814.640000 ;
      RECT 570.560000 814.010000 601.825000 814.640000 ;
      RECT 538.870000 814.010000 570.140000 814.640000 ;
      RECT 507.185000 814.010000 538.450000 814.640000 ;
      RECT 475.500000 814.010000 506.765000 814.640000 ;
      RECT 443.815000 814.010000 475.080000 814.640000 ;
      RECT 412.130000 814.010000 443.395000 814.640000 ;
      RECT 380.440000 814.010000 411.710000 814.640000 ;
      RECT 348.755000 814.010000 380.020000 814.640000 ;
      RECT 317.070000 814.010000 348.335000 814.640000 ;
      RECT 285.385000 814.010000 316.650000 814.640000 ;
      RECT 253.700000 814.010000 284.965000 814.640000 ;
      RECT 222.010000 814.010000 253.280000 814.640000 ;
      RECT 190.325000 814.010000 221.590000 814.640000 ;
      RECT 158.640000 814.010000 189.905000 814.640000 ;
      RECT 126.955000 814.010000 158.220000 814.640000 ;
      RECT 95.270000 814.010000 126.535000 814.640000 ;
      RECT 63.580000 814.010000 94.850000 814.640000 ;
      RECT 31.895000 814.010000 63.160000 814.640000 ;
      RECT 10.560000 814.010000 31.475000 814.640000 ;
      RECT 0.000000 814.010000 10.140000 814.015000 ;
      RECT 0.000000 0.630000 823.860000 814.010000 ;
      RECT 822.460000 0.000000 823.860000 0.630000 ;
      RECT 822.000000 0.000000 822.040000 0.630000 ;
      RECT 820.320000 0.000000 821.580000 0.630000 ;
      RECT 818.635000 0.000000 819.900000 0.630000 ;
      RECT 816.950000 0.000000 818.215000 0.630000 ;
      RECT 815.265000 0.000000 816.530000 0.630000 ;
      RECT 813.580000 0.000000 814.845000 0.630000 ;
      RECT 811.900000 0.000000 813.160000 0.630000 ;
      RECT 810.215000 0.000000 811.480000 0.630000 ;
      RECT 808.530000 0.000000 809.795000 0.630000 ;
      RECT 806.845000 0.000000 808.110000 0.630000 ;
      RECT 805.160000 0.000000 806.425000 0.630000 ;
      RECT 803.480000 0.000000 804.740000 0.630000 ;
      RECT 801.795000 0.000000 803.060000 0.630000 ;
      RECT 800.110000 0.000000 801.375000 0.630000 ;
      RECT 798.425000 0.000000 799.690000 0.630000 ;
      RECT 796.740000 0.000000 798.005000 0.630000 ;
      RECT 795.060000 0.000000 796.320000 0.630000 ;
      RECT 793.375000 0.000000 794.640000 0.630000 ;
      RECT 791.690000 0.000000 792.955000 0.630000 ;
      RECT 790.005000 0.000000 791.270000 0.630000 ;
      RECT 788.320000 0.000000 789.585000 0.630000 ;
      RECT 786.640000 0.000000 787.900000 0.630000 ;
      RECT 784.955000 0.000000 786.220000 0.630000 ;
      RECT 783.270000 0.000000 784.535000 0.630000 ;
      RECT 781.585000 0.000000 782.850000 0.630000 ;
      RECT 779.900000 0.000000 781.165000 0.630000 ;
      RECT 778.220000 0.000000 779.480000 0.630000 ;
      RECT 776.535000 0.000000 777.800000 0.630000 ;
      RECT 774.850000 0.000000 776.115000 0.630000 ;
      RECT 773.165000 0.000000 774.430000 0.630000 ;
      RECT 771.480000 0.000000 772.745000 0.630000 ;
      RECT 769.800000 0.000000 771.060000 0.630000 ;
      RECT 768.115000 0.000000 769.380000 0.630000 ;
      RECT 766.430000 0.000000 767.695000 0.630000 ;
      RECT 764.745000 0.000000 766.010000 0.630000 ;
      RECT 763.060000 0.000000 764.325000 0.630000 ;
      RECT 761.380000 0.000000 762.640000 0.630000 ;
      RECT 759.695000 0.000000 760.960000 0.630000 ;
      RECT 758.010000 0.000000 759.275000 0.630000 ;
      RECT 756.325000 0.000000 757.590000 0.630000 ;
      RECT 754.640000 0.000000 755.905000 0.630000 ;
      RECT 752.960000 0.000000 754.220000 0.630000 ;
      RECT 751.275000 0.000000 752.540000 0.630000 ;
      RECT 749.590000 0.000000 750.855000 0.630000 ;
      RECT 747.905000 0.000000 749.170000 0.630000 ;
      RECT 746.220000 0.000000 747.485000 0.630000 ;
      RECT 744.540000 0.000000 745.800000 0.630000 ;
      RECT 742.855000 0.000000 744.120000 0.630000 ;
      RECT 741.170000 0.000000 742.435000 0.630000 ;
      RECT 739.485000 0.000000 740.750000 0.630000 ;
      RECT 737.800000 0.000000 739.065000 0.630000 ;
      RECT 736.120000 0.000000 737.380000 0.630000 ;
      RECT 734.435000 0.000000 735.700000 0.630000 ;
      RECT 732.750000 0.000000 734.015000 0.630000 ;
      RECT 731.065000 0.000000 732.330000 0.630000 ;
      RECT 729.380000 0.000000 730.645000 0.630000 ;
      RECT 727.700000 0.000000 728.960000 0.630000 ;
      RECT 726.015000 0.000000 727.280000 0.630000 ;
      RECT 724.330000 0.000000 725.595000 0.630000 ;
      RECT 722.645000 0.000000 723.910000 0.630000 ;
      RECT 720.960000 0.000000 722.225000 0.630000 ;
      RECT 719.280000 0.000000 720.540000 0.630000 ;
      RECT 717.595000 0.000000 718.860000 0.630000 ;
      RECT 715.910000 0.000000 717.175000 0.630000 ;
      RECT 714.225000 0.000000 715.490000 0.630000 ;
      RECT 712.540000 0.000000 713.805000 0.630000 ;
      RECT 710.860000 0.000000 712.120000 0.630000 ;
      RECT 709.175000 0.000000 710.440000 0.630000 ;
      RECT 707.490000 0.000000 708.755000 0.630000 ;
      RECT 705.805000 0.000000 707.070000 0.630000 ;
      RECT 704.120000 0.000000 705.385000 0.630000 ;
      RECT 702.440000 0.000000 703.700000 0.630000 ;
      RECT 700.755000 0.000000 702.020000 0.630000 ;
      RECT 699.070000 0.000000 700.335000 0.630000 ;
      RECT 697.385000 0.000000 698.650000 0.630000 ;
      RECT 695.700000 0.000000 696.965000 0.630000 ;
      RECT 694.020000 0.000000 695.280000 0.630000 ;
      RECT 692.335000 0.000000 693.600000 0.630000 ;
      RECT 690.650000 0.000000 691.915000 0.630000 ;
      RECT 688.965000 0.000000 690.230000 0.630000 ;
      RECT 687.280000 0.000000 688.545000 0.630000 ;
      RECT 685.600000 0.000000 686.860000 0.630000 ;
      RECT 683.915000 0.000000 685.180000 0.630000 ;
      RECT 682.230000 0.000000 683.495000 0.630000 ;
      RECT 680.545000 0.000000 681.810000 0.630000 ;
      RECT 678.860000 0.000000 680.125000 0.630000 ;
      RECT 677.180000 0.000000 678.440000 0.630000 ;
      RECT 675.495000 0.000000 676.760000 0.630000 ;
      RECT 673.810000 0.000000 675.075000 0.630000 ;
      RECT 672.125000 0.000000 673.390000 0.630000 ;
      RECT 670.440000 0.000000 671.705000 0.630000 ;
      RECT 668.760000 0.000000 670.020000 0.630000 ;
      RECT 667.075000 0.000000 668.340000 0.630000 ;
      RECT 665.390000 0.000000 666.655000 0.630000 ;
      RECT 663.705000 0.000000 664.970000 0.630000 ;
      RECT 662.020000 0.000000 663.285000 0.630000 ;
      RECT 660.340000 0.000000 661.600000 0.630000 ;
      RECT 658.655000 0.000000 659.920000 0.630000 ;
      RECT 656.970000 0.000000 658.235000 0.630000 ;
      RECT 655.285000 0.000000 656.550000 0.630000 ;
      RECT 653.600000 0.000000 654.865000 0.630000 ;
      RECT 651.920000 0.000000 653.180000 0.630000 ;
      RECT 650.235000 0.000000 651.500000 0.630000 ;
      RECT 648.550000 0.000000 649.815000 0.630000 ;
      RECT 646.865000 0.000000 648.130000 0.630000 ;
      RECT 645.180000 0.000000 646.445000 0.630000 ;
      RECT 643.500000 0.000000 644.760000 0.630000 ;
      RECT 641.815000 0.000000 643.080000 0.630000 ;
      RECT 640.130000 0.000000 641.395000 0.630000 ;
      RECT 638.445000 0.000000 639.710000 0.630000 ;
      RECT 636.760000 0.000000 638.025000 0.630000 ;
      RECT 635.080000 0.000000 636.340000 0.630000 ;
      RECT 633.395000 0.000000 634.660000 0.630000 ;
      RECT 631.710000 0.000000 632.975000 0.630000 ;
      RECT 630.025000 0.000000 631.290000 0.630000 ;
      RECT 628.340000 0.000000 629.605000 0.630000 ;
      RECT 626.660000 0.000000 627.920000 0.630000 ;
      RECT 624.975000 0.000000 626.240000 0.630000 ;
      RECT 623.290000 0.000000 624.555000 0.630000 ;
      RECT 621.605000 0.000000 622.870000 0.630000 ;
      RECT 619.920000 0.000000 621.185000 0.630000 ;
      RECT 618.240000 0.000000 619.500000 0.630000 ;
      RECT 616.555000 0.000000 617.820000 0.630000 ;
      RECT 614.870000 0.000000 616.135000 0.630000 ;
      RECT 613.185000 0.000000 614.450000 0.630000 ;
      RECT 611.500000 0.000000 612.765000 0.630000 ;
      RECT 609.820000 0.000000 611.080000 0.630000 ;
      RECT 608.135000 0.000000 609.400000 0.630000 ;
      RECT 606.450000 0.000000 607.715000 0.630000 ;
      RECT 604.765000 0.000000 606.030000 0.630000 ;
      RECT 603.080000 0.000000 604.345000 0.630000 ;
      RECT 601.400000 0.000000 602.660000 0.630000 ;
      RECT 599.715000 0.000000 600.980000 0.630000 ;
      RECT 598.030000 0.000000 599.295000 0.630000 ;
      RECT 596.345000 0.000000 597.610000 0.630000 ;
      RECT 594.660000 0.000000 595.925000 0.630000 ;
      RECT 592.980000 0.000000 594.240000 0.630000 ;
      RECT 591.295000 0.000000 592.560000 0.630000 ;
      RECT 589.610000 0.000000 590.875000 0.630000 ;
      RECT 587.925000 0.000000 589.190000 0.630000 ;
      RECT 586.240000 0.000000 587.505000 0.630000 ;
      RECT 584.560000 0.000000 585.820000 0.630000 ;
      RECT 582.875000 0.000000 584.140000 0.630000 ;
      RECT 581.190000 0.000000 582.455000 0.630000 ;
      RECT 579.505000 0.000000 580.770000 0.630000 ;
      RECT 577.820000 0.000000 579.085000 0.630000 ;
      RECT 576.140000 0.000000 577.400000 0.630000 ;
      RECT 574.455000 0.000000 575.720000 0.630000 ;
      RECT 572.770000 0.000000 574.035000 0.630000 ;
      RECT 571.085000 0.000000 572.350000 0.630000 ;
      RECT 569.400000 0.000000 570.665000 0.630000 ;
      RECT 567.720000 0.000000 568.980000 0.630000 ;
      RECT 566.035000 0.000000 567.300000 0.630000 ;
      RECT 564.350000 0.000000 565.615000 0.630000 ;
      RECT 562.665000 0.000000 563.930000 0.630000 ;
      RECT 560.980000 0.000000 562.245000 0.630000 ;
      RECT 559.300000 0.000000 560.560000 0.630000 ;
      RECT 557.615000 0.000000 558.880000 0.630000 ;
      RECT 555.930000 0.000000 557.195000 0.630000 ;
      RECT 554.245000 0.000000 555.510000 0.630000 ;
      RECT 552.560000 0.000000 553.825000 0.630000 ;
      RECT 550.880000 0.000000 552.140000 0.630000 ;
      RECT 549.195000 0.000000 550.460000 0.630000 ;
      RECT 547.510000 0.000000 548.775000 0.630000 ;
      RECT 545.825000 0.000000 547.090000 0.630000 ;
      RECT 544.140000 0.000000 545.405000 0.630000 ;
      RECT 542.460000 0.000000 543.720000 0.630000 ;
      RECT 540.775000 0.000000 542.040000 0.630000 ;
      RECT 539.090000 0.000000 540.355000 0.630000 ;
      RECT 537.405000 0.000000 538.670000 0.630000 ;
      RECT 535.720000 0.000000 536.985000 0.630000 ;
      RECT 534.040000 0.000000 535.300000 0.630000 ;
      RECT 532.355000 0.000000 533.620000 0.630000 ;
      RECT 530.670000 0.000000 531.935000 0.630000 ;
      RECT 528.985000 0.000000 530.250000 0.630000 ;
      RECT 527.300000 0.000000 528.565000 0.630000 ;
      RECT 525.620000 0.000000 526.880000 0.630000 ;
      RECT 523.935000 0.000000 525.200000 0.630000 ;
      RECT 522.250000 0.000000 523.515000 0.630000 ;
      RECT 520.565000 0.000000 521.830000 0.630000 ;
      RECT 518.880000 0.000000 520.145000 0.630000 ;
      RECT 517.200000 0.000000 518.460000 0.630000 ;
      RECT 515.515000 0.000000 516.780000 0.630000 ;
      RECT 513.830000 0.000000 515.095000 0.630000 ;
      RECT 512.145000 0.000000 513.410000 0.630000 ;
      RECT 510.460000 0.000000 511.725000 0.630000 ;
      RECT 508.780000 0.000000 510.040000 0.630000 ;
      RECT 507.095000 0.000000 508.360000 0.630000 ;
      RECT 505.410000 0.000000 506.675000 0.630000 ;
      RECT 503.725000 0.000000 504.990000 0.630000 ;
      RECT 502.040000 0.000000 503.305000 0.630000 ;
      RECT 500.360000 0.000000 501.620000 0.630000 ;
      RECT 498.675000 0.000000 499.940000 0.630000 ;
      RECT 496.990000 0.000000 498.255000 0.630000 ;
      RECT 495.305000 0.000000 496.570000 0.630000 ;
      RECT 493.620000 0.000000 494.885000 0.630000 ;
      RECT 491.940000 0.000000 493.200000 0.630000 ;
      RECT 490.255000 0.000000 491.520000 0.630000 ;
      RECT 488.570000 0.000000 489.835000 0.630000 ;
      RECT 486.885000 0.000000 488.150000 0.630000 ;
      RECT 485.200000 0.000000 486.465000 0.630000 ;
      RECT 483.520000 0.000000 484.780000 0.630000 ;
      RECT 481.835000 0.000000 483.100000 0.630000 ;
      RECT 480.150000 0.000000 481.415000 0.630000 ;
      RECT 478.465000 0.000000 479.730000 0.630000 ;
      RECT 476.780000 0.000000 478.045000 0.630000 ;
      RECT 475.100000 0.000000 476.360000 0.630000 ;
      RECT 473.415000 0.000000 474.680000 0.630000 ;
      RECT 471.730000 0.000000 472.995000 0.630000 ;
      RECT 470.045000 0.000000 471.310000 0.630000 ;
      RECT 468.360000 0.000000 469.625000 0.630000 ;
      RECT 466.680000 0.000000 467.940000 0.630000 ;
      RECT 464.995000 0.000000 466.260000 0.630000 ;
      RECT 463.310000 0.000000 464.575000 0.630000 ;
      RECT 461.625000 0.000000 462.890000 0.630000 ;
      RECT 459.940000 0.000000 461.205000 0.630000 ;
      RECT 458.260000 0.000000 459.520000 0.630000 ;
      RECT 456.575000 0.000000 457.840000 0.630000 ;
      RECT 454.890000 0.000000 456.155000 0.630000 ;
      RECT 453.205000 0.000000 454.470000 0.630000 ;
      RECT 451.520000 0.000000 452.785000 0.630000 ;
      RECT 449.840000 0.000000 451.100000 0.630000 ;
      RECT 448.155000 0.000000 449.420000 0.630000 ;
      RECT 446.470000 0.000000 447.735000 0.630000 ;
      RECT 444.785000 0.000000 446.050000 0.630000 ;
      RECT 443.100000 0.000000 444.365000 0.630000 ;
      RECT 441.420000 0.000000 442.680000 0.630000 ;
      RECT 439.735000 0.000000 441.000000 0.630000 ;
      RECT 438.050000 0.000000 439.315000 0.630000 ;
      RECT 436.365000 0.000000 437.630000 0.630000 ;
      RECT 434.680000 0.000000 435.945000 0.630000 ;
      RECT 433.000000 0.000000 434.260000 0.630000 ;
      RECT 431.315000 0.000000 432.580000 0.630000 ;
      RECT 429.630000 0.000000 430.895000 0.630000 ;
      RECT 427.945000 0.000000 429.210000 0.630000 ;
      RECT 426.260000 0.000000 427.525000 0.630000 ;
      RECT 424.580000 0.000000 425.840000 0.630000 ;
      RECT 422.895000 0.000000 424.160000 0.630000 ;
      RECT 421.210000 0.000000 422.475000 0.630000 ;
      RECT 419.525000 0.000000 420.790000 0.630000 ;
      RECT 417.840000 0.000000 419.105000 0.630000 ;
      RECT 416.160000 0.000000 417.420000 0.630000 ;
      RECT 414.475000 0.000000 415.740000 0.630000 ;
      RECT 412.790000 0.000000 414.055000 0.630000 ;
      RECT 411.105000 0.000000 412.370000 0.630000 ;
      RECT 409.420000 0.000000 410.685000 0.630000 ;
      RECT 407.740000 0.000000 409.000000 0.630000 ;
      RECT 406.055000 0.000000 407.320000 0.630000 ;
      RECT 404.370000 0.000000 405.635000 0.630000 ;
      RECT 402.685000 0.000000 403.950000 0.630000 ;
      RECT 401.000000 0.000000 402.265000 0.630000 ;
      RECT 399.320000 0.000000 400.580000 0.630000 ;
      RECT 397.635000 0.000000 398.900000 0.630000 ;
      RECT 395.950000 0.000000 397.215000 0.630000 ;
      RECT 394.265000 0.000000 395.530000 0.630000 ;
      RECT 392.580000 0.000000 393.845000 0.630000 ;
      RECT 390.900000 0.000000 392.160000 0.630000 ;
      RECT 389.215000 0.000000 390.480000 0.630000 ;
      RECT 387.530000 0.000000 388.795000 0.630000 ;
      RECT 385.845000 0.000000 387.110000 0.630000 ;
      RECT 384.160000 0.000000 385.425000 0.630000 ;
      RECT 382.480000 0.000000 383.740000 0.630000 ;
      RECT 380.795000 0.000000 382.060000 0.630000 ;
      RECT 379.110000 0.000000 380.375000 0.630000 ;
      RECT 377.425000 0.000000 378.690000 0.630000 ;
      RECT 375.740000 0.000000 377.005000 0.630000 ;
      RECT 374.060000 0.000000 375.320000 0.630000 ;
      RECT 372.375000 0.000000 373.640000 0.630000 ;
      RECT 370.690000 0.000000 371.955000 0.630000 ;
      RECT 369.005000 0.000000 370.270000 0.630000 ;
      RECT 367.320000 0.000000 368.585000 0.630000 ;
      RECT 365.640000 0.000000 366.900000 0.630000 ;
      RECT 363.955000 0.000000 365.220000 0.630000 ;
      RECT 362.270000 0.000000 363.535000 0.630000 ;
      RECT 360.585000 0.000000 361.850000 0.630000 ;
      RECT 358.900000 0.000000 360.165000 0.630000 ;
      RECT 357.220000 0.000000 358.480000 0.630000 ;
      RECT 355.535000 0.000000 356.800000 0.630000 ;
      RECT 353.850000 0.000000 355.115000 0.630000 ;
      RECT 352.165000 0.000000 353.430000 0.630000 ;
      RECT 350.480000 0.000000 351.745000 0.630000 ;
      RECT 348.800000 0.000000 350.060000 0.630000 ;
      RECT 347.115000 0.000000 348.380000 0.630000 ;
      RECT 345.430000 0.000000 346.695000 0.630000 ;
      RECT 343.745000 0.000000 345.010000 0.630000 ;
      RECT 342.060000 0.000000 343.325000 0.630000 ;
      RECT 340.380000 0.000000 341.640000 0.630000 ;
      RECT 338.695000 0.000000 339.960000 0.630000 ;
      RECT 337.010000 0.000000 338.275000 0.630000 ;
      RECT 335.325000 0.000000 336.590000 0.630000 ;
      RECT 333.640000 0.000000 334.905000 0.630000 ;
      RECT 331.960000 0.000000 333.220000 0.630000 ;
      RECT 330.275000 0.000000 331.540000 0.630000 ;
      RECT 328.590000 0.000000 329.855000 0.630000 ;
      RECT 326.905000 0.000000 328.170000 0.630000 ;
      RECT 325.220000 0.000000 326.485000 0.630000 ;
      RECT 323.540000 0.000000 324.800000 0.630000 ;
      RECT 321.855000 0.000000 323.120000 0.630000 ;
      RECT 320.170000 0.000000 321.435000 0.630000 ;
      RECT 318.485000 0.000000 319.750000 0.630000 ;
      RECT 316.800000 0.000000 318.065000 0.630000 ;
      RECT 315.120000 0.000000 316.380000 0.630000 ;
      RECT 313.435000 0.000000 314.700000 0.630000 ;
      RECT 311.750000 0.000000 313.015000 0.630000 ;
      RECT 310.065000 0.000000 311.330000 0.630000 ;
      RECT 308.380000 0.000000 309.645000 0.630000 ;
      RECT 306.700000 0.000000 307.960000 0.630000 ;
      RECT 305.015000 0.000000 306.280000 0.630000 ;
      RECT 303.330000 0.000000 304.595000 0.630000 ;
      RECT 301.645000 0.000000 302.910000 0.630000 ;
      RECT 299.960000 0.000000 301.225000 0.630000 ;
      RECT 298.280000 0.000000 299.540000 0.630000 ;
      RECT 296.595000 0.000000 297.860000 0.630000 ;
      RECT 294.910000 0.000000 296.175000 0.630000 ;
      RECT 293.225000 0.000000 294.490000 0.630000 ;
      RECT 291.540000 0.000000 292.805000 0.630000 ;
      RECT 289.860000 0.000000 291.120000 0.630000 ;
      RECT 288.175000 0.000000 289.440000 0.630000 ;
      RECT 286.490000 0.000000 287.755000 0.630000 ;
      RECT 284.805000 0.000000 286.070000 0.630000 ;
      RECT 283.120000 0.000000 284.385000 0.630000 ;
      RECT 281.440000 0.000000 282.700000 0.630000 ;
      RECT 279.755000 0.000000 281.020000 0.630000 ;
      RECT 278.070000 0.000000 279.335000 0.630000 ;
      RECT 276.385000 0.000000 277.650000 0.630000 ;
      RECT 274.700000 0.000000 275.965000 0.630000 ;
      RECT 273.020000 0.000000 274.280000 0.630000 ;
      RECT 271.335000 0.000000 272.600000 0.630000 ;
      RECT 269.650000 0.000000 270.915000 0.630000 ;
      RECT 267.965000 0.000000 269.230000 0.630000 ;
      RECT 266.280000 0.000000 267.545000 0.630000 ;
      RECT 264.600000 0.000000 265.860000 0.630000 ;
      RECT 262.915000 0.000000 264.180000 0.630000 ;
      RECT 261.230000 0.000000 262.495000 0.630000 ;
      RECT 259.545000 0.000000 260.810000 0.630000 ;
      RECT 257.860000 0.000000 259.125000 0.630000 ;
      RECT 256.180000 0.000000 257.440000 0.630000 ;
      RECT 254.495000 0.000000 255.760000 0.630000 ;
      RECT 252.810000 0.000000 254.075000 0.630000 ;
      RECT 251.125000 0.000000 252.390000 0.630000 ;
      RECT 249.440000 0.000000 250.705000 0.630000 ;
      RECT 247.760000 0.000000 249.020000 0.630000 ;
      RECT 246.075000 0.000000 247.340000 0.630000 ;
      RECT 244.390000 0.000000 245.655000 0.630000 ;
      RECT 242.705000 0.000000 243.970000 0.630000 ;
      RECT 241.020000 0.000000 242.285000 0.630000 ;
      RECT 239.340000 0.000000 240.600000 0.630000 ;
      RECT 237.655000 0.000000 238.920000 0.630000 ;
      RECT 235.970000 0.000000 237.235000 0.630000 ;
      RECT 234.285000 0.000000 235.550000 0.630000 ;
      RECT 232.600000 0.000000 233.865000 0.630000 ;
      RECT 230.920000 0.000000 232.180000 0.630000 ;
      RECT 229.235000 0.000000 230.500000 0.630000 ;
      RECT 227.550000 0.000000 228.815000 0.630000 ;
      RECT 225.865000 0.000000 227.130000 0.630000 ;
      RECT 224.180000 0.000000 225.445000 0.630000 ;
      RECT 222.500000 0.000000 223.760000 0.630000 ;
      RECT 220.815000 0.000000 222.080000 0.630000 ;
      RECT 219.130000 0.000000 220.395000 0.630000 ;
      RECT 217.445000 0.000000 218.710000 0.630000 ;
      RECT 215.760000 0.000000 217.025000 0.630000 ;
      RECT 214.080000 0.000000 215.340000 0.630000 ;
      RECT 212.395000 0.000000 213.660000 0.630000 ;
      RECT 210.710000 0.000000 211.975000 0.630000 ;
      RECT 209.025000 0.000000 210.290000 0.630000 ;
      RECT 207.340000 0.000000 208.605000 0.630000 ;
      RECT 205.660000 0.000000 206.920000 0.630000 ;
      RECT 203.975000 0.000000 205.240000 0.630000 ;
      RECT 202.290000 0.000000 203.555000 0.630000 ;
      RECT 200.605000 0.000000 201.870000 0.630000 ;
      RECT 198.920000 0.000000 200.185000 0.630000 ;
      RECT 197.240000 0.000000 198.500000 0.630000 ;
      RECT 195.555000 0.000000 196.820000 0.630000 ;
      RECT 193.870000 0.000000 195.135000 0.630000 ;
      RECT 192.185000 0.000000 193.450000 0.630000 ;
      RECT 190.500000 0.000000 191.765000 0.630000 ;
      RECT 188.820000 0.000000 190.080000 0.630000 ;
      RECT 187.135000 0.000000 188.400000 0.630000 ;
      RECT 185.450000 0.000000 186.715000 0.630000 ;
      RECT 183.765000 0.000000 185.030000 0.630000 ;
      RECT 182.080000 0.000000 183.345000 0.630000 ;
      RECT 180.400000 0.000000 181.660000 0.630000 ;
      RECT 178.715000 0.000000 179.980000 0.630000 ;
      RECT 177.030000 0.000000 178.295000 0.630000 ;
      RECT 175.345000 0.000000 176.610000 0.630000 ;
      RECT 173.660000 0.000000 174.925000 0.630000 ;
      RECT 171.980000 0.000000 173.240000 0.630000 ;
      RECT 170.295000 0.000000 171.560000 0.630000 ;
      RECT 168.610000 0.000000 169.875000 0.630000 ;
      RECT 166.925000 0.000000 168.190000 0.630000 ;
      RECT 165.240000 0.000000 166.505000 0.630000 ;
      RECT 163.560000 0.000000 164.820000 0.630000 ;
      RECT 161.875000 0.000000 163.140000 0.630000 ;
      RECT 160.190000 0.000000 161.455000 0.630000 ;
      RECT 158.505000 0.000000 159.770000 0.630000 ;
      RECT 156.820000 0.000000 158.085000 0.630000 ;
      RECT 155.140000 0.000000 156.400000 0.630000 ;
      RECT 153.455000 0.000000 154.720000 0.630000 ;
      RECT 151.770000 0.000000 153.035000 0.630000 ;
      RECT 150.085000 0.000000 151.350000 0.630000 ;
      RECT 148.400000 0.000000 149.665000 0.630000 ;
      RECT 146.720000 0.000000 147.980000 0.630000 ;
      RECT 145.035000 0.000000 146.300000 0.630000 ;
      RECT 143.350000 0.000000 144.615000 0.630000 ;
      RECT 141.665000 0.000000 142.930000 0.630000 ;
      RECT 139.980000 0.000000 141.245000 0.630000 ;
      RECT 138.300000 0.000000 139.560000 0.630000 ;
      RECT 136.615000 0.000000 137.880000 0.630000 ;
      RECT 134.930000 0.000000 136.195000 0.630000 ;
      RECT 133.245000 0.000000 134.510000 0.630000 ;
      RECT 131.560000 0.000000 132.825000 0.630000 ;
      RECT 129.880000 0.000000 131.140000 0.630000 ;
      RECT 128.195000 0.000000 129.460000 0.630000 ;
      RECT 126.510000 0.000000 127.775000 0.630000 ;
      RECT 124.825000 0.000000 126.090000 0.630000 ;
      RECT 123.140000 0.000000 124.405000 0.630000 ;
      RECT 121.460000 0.000000 122.720000 0.630000 ;
      RECT 119.775000 0.000000 121.040000 0.630000 ;
      RECT 118.090000 0.000000 119.355000 0.630000 ;
      RECT 116.405000 0.000000 117.670000 0.630000 ;
      RECT 114.720000 0.000000 115.985000 0.630000 ;
      RECT 113.040000 0.000000 114.300000 0.630000 ;
      RECT 111.355000 0.000000 112.620000 0.630000 ;
      RECT 109.670000 0.000000 110.935000 0.630000 ;
      RECT 107.985000 0.000000 109.250000 0.630000 ;
      RECT 106.300000 0.000000 107.565000 0.630000 ;
      RECT 104.620000 0.000000 105.880000 0.630000 ;
      RECT 102.935000 0.000000 104.200000 0.630000 ;
      RECT 101.250000 0.000000 102.515000 0.630000 ;
      RECT 99.565000 0.000000 100.830000 0.630000 ;
      RECT 97.880000 0.000000 99.145000 0.630000 ;
      RECT 96.200000 0.000000 97.460000 0.630000 ;
      RECT 94.515000 0.000000 95.780000 0.630000 ;
      RECT 92.830000 0.000000 94.095000 0.630000 ;
      RECT 91.145000 0.000000 92.410000 0.630000 ;
      RECT 89.460000 0.000000 90.725000 0.630000 ;
      RECT 87.780000 0.000000 89.040000 0.630000 ;
      RECT 86.095000 0.000000 87.360000 0.630000 ;
      RECT 84.410000 0.000000 85.675000 0.630000 ;
      RECT 82.725000 0.000000 83.990000 0.630000 ;
      RECT 81.040000 0.000000 82.305000 0.630000 ;
      RECT 79.360000 0.000000 80.620000 0.630000 ;
      RECT 77.675000 0.000000 78.940000 0.630000 ;
      RECT 75.990000 0.000000 77.255000 0.630000 ;
      RECT 74.305000 0.000000 75.570000 0.630000 ;
      RECT 72.620000 0.000000 73.885000 0.630000 ;
      RECT 70.940000 0.000000 72.200000 0.630000 ;
      RECT 69.255000 0.000000 70.520000 0.630000 ;
      RECT 67.570000 0.000000 68.835000 0.630000 ;
      RECT 65.885000 0.000000 67.150000 0.630000 ;
      RECT 64.200000 0.000000 65.465000 0.630000 ;
      RECT 62.520000 0.000000 63.780000 0.630000 ;
      RECT 60.835000 0.000000 62.100000 0.630000 ;
      RECT 59.150000 0.000000 60.415000 0.630000 ;
      RECT 57.465000 0.000000 58.730000 0.630000 ;
      RECT 55.780000 0.000000 57.045000 0.630000 ;
      RECT 54.100000 0.000000 55.360000 0.630000 ;
      RECT 52.415000 0.000000 53.680000 0.630000 ;
      RECT 50.730000 0.000000 51.995000 0.630000 ;
      RECT 49.045000 0.000000 50.310000 0.630000 ;
      RECT 47.360000 0.000000 48.625000 0.630000 ;
      RECT 45.680000 0.000000 46.940000 0.630000 ;
      RECT 43.995000 0.000000 45.260000 0.630000 ;
      RECT 42.310000 0.000000 43.575000 0.630000 ;
      RECT 40.625000 0.000000 41.890000 0.630000 ;
      RECT 38.940000 0.000000 40.205000 0.630000 ;
      RECT 37.260000 0.000000 38.520000 0.630000 ;
      RECT 35.575000 0.000000 36.840000 0.630000 ;
      RECT 33.890000 0.000000 35.155000 0.630000 ;
      RECT 32.205000 0.000000 33.470000 0.630000 ;
      RECT 30.520000 0.000000 31.785000 0.630000 ;
      RECT 28.840000 0.000000 30.100000 0.630000 ;
      RECT 27.155000 0.000000 28.420000 0.630000 ;
      RECT 25.470000 0.000000 26.735000 0.630000 ;
      RECT 23.785000 0.000000 25.050000 0.630000 ;
      RECT 22.100000 0.000000 23.365000 0.630000 ;
      RECT 20.420000 0.000000 21.680000 0.630000 ;
      RECT 18.735000 0.000000 20.000000 0.630000 ;
      RECT 17.050000 0.000000 18.315000 0.630000 ;
      RECT 15.365000 0.000000 16.630000 0.630000 ;
      RECT 13.680000 0.000000 14.945000 0.630000 ;
      RECT 12.000000 0.000000 13.260000 0.630000 ;
      RECT 10.315000 0.000000 11.580000 0.630000 ;
      RECT 8.630000 0.000000 9.895000 0.630000 ;
      RECT 6.945000 0.000000 8.210000 0.630000 ;
      RECT 5.260000 0.000000 6.525000 0.630000 ;
      RECT 3.580000 0.000000 4.840000 0.630000 ;
      RECT 1.895000 0.000000 3.160000 0.630000 ;
      RECT 0.900000 0.000000 1.475000 0.630000 ;
      RECT 0.000000 0.000000 0.480000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 811.140000 823.860000 814.640000 ;
      RECT 1.100000 810.530000 823.860000 811.140000 ;
      RECT 1.100000 810.240000 822.760000 810.530000 ;
      RECT 0.000000 809.630000 822.760000 810.240000 ;
      RECT 0.000000 796.550000 823.860000 809.630000 ;
      RECT 0.000000 795.650000 822.760000 796.550000 ;
      RECT 0.000000 795.210000 823.860000 795.650000 ;
      RECT 1.100000 794.310000 823.860000 795.210000 ;
      RECT 0.000000 778.040000 823.860000 794.310000 ;
      RECT 0.000000 777.140000 822.760000 778.040000 ;
      RECT 0.000000 775.340000 823.860000 777.140000 ;
      RECT 1.100000 774.440000 823.860000 775.340000 ;
      RECT 0.000000 759.525000 823.860000 774.440000 ;
      RECT 0.000000 758.625000 822.760000 759.525000 ;
      RECT 0.000000 755.470000 823.860000 758.625000 ;
      RECT 1.100000 754.570000 823.860000 755.470000 ;
      RECT 0.000000 741.010000 823.860000 754.570000 ;
      RECT 0.000000 740.110000 822.760000 741.010000 ;
      RECT 0.000000 735.605000 823.860000 740.110000 ;
      RECT 1.100000 734.705000 823.860000 735.605000 ;
      RECT 0.000000 722.495000 823.860000 734.705000 ;
      RECT 0.000000 721.595000 822.760000 722.495000 ;
      RECT 0.000000 715.735000 823.860000 721.595000 ;
      RECT 1.100000 714.835000 823.860000 715.735000 ;
      RECT 0.000000 703.980000 823.860000 714.835000 ;
      RECT 0.000000 703.080000 822.760000 703.980000 ;
      RECT 0.000000 695.865000 823.860000 703.080000 ;
      RECT 1.100000 694.965000 823.860000 695.865000 ;
      RECT 0.000000 685.470000 823.860000 694.965000 ;
      RECT 0.000000 684.570000 822.760000 685.470000 ;
      RECT 0.000000 675.995000 823.860000 684.570000 ;
      RECT 1.100000 675.095000 823.860000 675.995000 ;
      RECT 0.000000 666.955000 823.860000 675.095000 ;
      RECT 0.000000 666.055000 822.760000 666.955000 ;
      RECT 0.000000 656.125000 823.860000 666.055000 ;
      RECT 1.100000 655.225000 823.860000 656.125000 ;
      RECT 0.000000 648.440000 823.860000 655.225000 ;
      RECT 0.000000 647.540000 822.760000 648.440000 ;
      RECT 0.000000 636.260000 823.860000 647.540000 ;
      RECT 1.100000 635.360000 823.860000 636.260000 ;
      RECT 0.000000 629.925000 823.860000 635.360000 ;
      RECT 0.000000 629.025000 822.760000 629.925000 ;
      RECT 0.000000 616.390000 823.860000 629.025000 ;
      RECT 1.100000 615.490000 823.860000 616.390000 ;
      RECT 0.000000 611.410000 823.860000 615.490000 ;
      RECT 0.000000 610.510000 822.760000 611.410000 ;
      RECT 0.000000 596.520000 823.860000 610.510000 ;
      RECT 1.100000 595.620000 823.860000 596.520000 ;
      RECT 0.000000 592.900000 823.860000 595.620000 ;
      RECT 0.000000 592.000000 822.760000 592.900000 ;
      RECT 0.000000 576.650000 823.860000 592.000000 ;
      RECT 1.100000 575.750000 823.860000 576.650000 ;
      RECT 0.000000 574.385000 823.860000 575.750000 ;
      RECT 0.000000 573.485000 822.760000 574.385000 ;
      RECT 0.000000 556.780000 823.860000 573.485000 ;
      RECT 1.100000 555.880000 823.860000 556.780000 ;
      RECT 0.000000 555.870000 823.860000 555.880000 ;
      RECT 0.000000 554.970000 822.760000 555.870000 ;
      RECT 0.000000 537.355000 823.860000 554.970000 ;
      RECT 0.000000 536.915000 822.760000 537.355000 ;
      RECT 1.100000 536.455000 822.760000 536.915000 ;
      RECT 1.100000 536.015000 823.860000 536.455000 ;
      RECT 0.000000 518.840000 823.860000 536.015000 ;
      RECT 0.000000 517.940000 822.760000 518.840000 ;
      RECT 0.000000 517.045000 823.860000 517.940000 ;
      RECT 1.100000 516.145000 823.860000 517.045000 ;
      RECT 0.000000 500.330000 823.860000 516.145000 ;
      RECT 0.000000 499.430000 822.760000 500.330000 ;
      RECT 0.000000 497.175000 823.860000 499.430000 ;
      RECT 1.100000 496.275000 823.860000 497.175000 ;
      RECT 0.000000 481.815000 823.860000 496.275000 ;
      RECT 0.000000 480.915000 822.760000 481.815000 ;
      RECT 0.000000 477.305000 823.860000 480.915000 ;
      RECT 1.100000 476.405000 823.860000 477.305000 ;
      RECT 0.000000 463.300000 823.860000 476.405000 ;
      RECT 0.000000 462.400000 822.760000 463.300000 ;
      RECT 0.000000 457.435000 823.860000 462.400000 ;
      RECT 1.100000 456.535000 823.860000 457.435000 ;
      RECT 0.000000 444.785000 823.860000 456.535000 ;
      RECT 0.000000 443.885000 822.760000 444.785000 ;
      RECT 0.000000 437.570000 823.860000 443.885000 ;
      RECT 1.100000 436.670000 823.860000 437.570000 ;
      RECT 0.000000 426.270000 823.860000 436.670000 ;
      RECT 0.000000 425.370000 822.760000 426.270000 ;
      RECT 0.000000 417.700000 823.860000 425.370000 ;
      RECT 1.100000 416.800000 823.860000 417.700000 ;
      RECT 0.000000 407.760000 823.860000 416.800000 ;
      RECT 0.000000 406.860000 822.760000 407.760000 ;
      RECT 0.000000 397.830000 823.860000 406.860000 ;
      RECT 1.100000 396.930000 823.860000 397.830000 ;
      RECT 0.000000 389.245000 823.860000 396.930000 ;
      RECT 0.000000 388.345000 822.760000 389.245000 ;
      RECT 0.000000 384.750000 823.860000 388.345000 ;
      RECT 0.000000 382.150000 821.560000 384.750000 ;
      RECT 0.000000 380.750000 823.860000 382.150000 ;
      RECT 0.000000 378.150000 821.560000 380.750000 ;
      RECT 0.000000 377.960000 823.860000 378.150000 ;
      RECT 1.100000 377.060000 823.860000 377.960000 ;
      RECT 0.000000 370.730000 823.860000 377.060000 ;
      RECT 0.000000 369.830000 822.760000 370.730000 ;
      RECT 0.000000 358.090000 823.860000 369.830000 ;
      RECT 1.100000 357.190000 823.860000 358.090000 ;
      RECT 0.000000 352.215000 823.860000 357.190000 ;
      RECT 0.000000 351.315000 822.760000 352.215000 ;
      RECT 0.000000 338.225000 823.860000 351.315000 ;
      RECT 1.100000 337.325000 823.860000 338.225000 ;
      RECT 0.000000 333.700000 823.860000 337.325000 ;
      RECT 0.000000 332.800000 822.760000 333.700000 ;
      RECT 0.000000 318.355000 823.860000 332.800000 ;
      RECT 1.100000 317.455000 823.860000 318.355000 ;
      RECT 0.000000 315.190000 823.860000 317.455000 ;
      RECT 0.000000 314.290000 822.760000 315.190000 ;
      RECT 0.000000 298.485000 823.860000 314.290000 ;
      RECT 1.100000 297.585000 823.860000 298.485000 ;
      RECT 0.000000 296.675000 823.860000 297.585000 ;
      RECT 0.000000 295.775000 822.760000 296.675000 ;
      RECT 0.000000 278.615000 823.860000 295.775000 ;
      RECT 1.100000 278.160000 823.860000 278.615000 ;
      RECT 1.100000 277.715000 822.760000 278.160000 ;
      RECT 0.000000 277.260000 822.760000 277.715000 ;
      RECT 0.000000 259.645000 823.860000 277.260000 ;
      RECT 0.000000 258.745000 822.760000 259.645000 ;
      RECT 1.100000 257.845000 823.860000 258.745000 ;
      RECT 0.000000 241.130000 823.860000 257.845000 ;
      RECT 0.000000 240.230000 822.760000 241.130000 ;
      RECT 0.000000 238.880000 823.860000 240.230000 ;
      RECT 1.100000 237.980000 823.860000 238.880000 ;
      RECT 0.000000 222.620000 823.860000 237.980000 ;
      RECT 0.000000 221.720000 822.760000 222.620000 ;
      RECT 0.000000 219.010000 823.860000 221.720000 ;
      RECT 1.100000 218.110000 823.860000 219.010000 ;
      RECT 0.000000 204.105000 823.860000 218.110000 ;
      RECT 0.000000 203.205000 822.760000 204.105000 ;
      RECT 0.000000 199.140000 823.860000 203.205000 ;
      RECT 1.100000 198.240000 823.860000 199.140000 ;
      RECT 0.000000 185.590000 823.860000 198.240000 ;
      RECT 0.000000 184.690000 822.760000 185.590000 ;
      RECT 0.000000 179.270000 823.860000 184.690000 ;
      RECT 1.100000 178.370000 823.860000 179.270000 ;
      RECT 0.000000 167.075000 823.860000 178.370000 ;
      RECT 0.000000 166.175000 822.760000 167.075000 ;
      RECT 0.000000 159.400000 823.860000 166.175000 ;
      RECT 1.100000 158.500000 823.860000 159.400000 ;
      RECT 0.000000 148.560000 823.860000 158.500000 ;
      RECT 0.000000 147.660000 822.760000 148.560000 ;
      RECT 0.000000 139.535000 823.860000 147.660000 ;
      RECT 1.100000 138.635000 823.860000 139.535000 ;
      RECT 0.000000 130.050000 823.860000 138.635000 ;
      RECT 0.000000 129.150000 822.760000 130.050000 ;
      RECT 0.000000 119.665000 823.860000 129.150000 ;
      RECT 1.100000 118.765000 823.860000 119.665000 ;
      RECT 0.000000 111.535000 823.860000 118.765000 ;
      RECT 0.000000 110.635000 822.760000 111.535000 ;
      RECT 0.000000 99.795000 823.860000 110.635000 ;
      RECT 1.100000 98.895000 823.860000 99.795000 ;
      RECT 0.000000 93.020000 823.860000 98.895000 ;
      RECT 0.000000 92.120000 822.760000 93.020000 ;
      RECT 0.000000 79.925000 823.860000 92.120000 ;
      RECT 1.100000 79.025000 823.860000 79.925000 ;
      RECT 0.000000 74.505000 823.860000 79.025000 ;
      RECT 0.000000 73.605000 822.760000 74.505000 ;
      RECT 0.000000 60.055000 823.860000 73.605000 ;
      RECT 1.100000 59.155000 823.860000 60.055000 ;
      RECT 0.000000 55.990000 823.860000 59.155000 ;
      RECT 0.000000 55.090000 822.760000 55.990000 ;
      RECT 0.000000 40.190000 823.860000 55.090000 ;
      RECT 1.100000 39.290000 823.860000 40.190000 ;
      RECT 0.000000 37.480000 823.860000 39.290000 ;
      RECT 0.000000 36.580000 822.760000 37.480000 ;
      RECT 0.000000 20.320000 823.860000 36.580000 ;
      RECT 1.100000 19.420000 823.860000 20.320000 ;
      RECT 0.000000 18.965000 823.860000 19.420000 ;
      RECT 0.000000 18.065000 822.760000 18.965000 ;
      RECT 0.000000 10.820000 823.860000 18.065000 ;
      RECT 1.100000 10.210000 823.860000 10.820000 ;
      RECT 1.100000 9.920000 822.760000 10.210000 ;
      RECT 0.000000 9.310000 822.760000 9.920000 ;
      RECT 0.000000 0.000000 823.860000 9.310000 ;
    LAYER met4 ;
      RECT 311.765000 812.840000 823.860000 814.640000 ;
      RECT 0.000000 812.840000 305.165000 814.640000 ;
      RECT 311.765000 812.340000 819.500000 812.840000 ;
      RECT 307.765000 812.340000 309.165000 814.640000 ;
      RECT 4.360000 812.340000 305.165000 812.840000 ;
      RECT 4.360000 808.840000 819.500000 812.340000 ;
      RECT 818.100000 5.800000 819.500000 808.840000 ;
      RECT 8.360000 5.800000 815.500000 808.840000 ;
      RECT 4.360000 5.800000 5.760000 808.840000 ;
      RECT 822.100000 1.800000 823.860000 812.840000 ;
      RECT 817.300000 1.800000 819.500000 5.800000 ;
      RECT 4.360000 1.800000 815.500000 5.800000 ;
      RECT 0.000000 1.800000 1.760000 812.840000 ;
      RECT 817.300000 0.500000 823.860000 1.800000 ;
      RECT 0.000000 0.500000 815.500000 1.800000 ;
      RECT 0.000000 0.000000 823.860000 0.500000 ;
  END
END user_proj_example

END LIBRARY
